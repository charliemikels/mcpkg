module mcpkg

fn platform_modrinth() ModPlatform {
	return ModPlatform {
		name: 'modrinth'
		home_url: 'https://modrinth.com/'
	}
}
