module mcpkg

struct BranchJson {}

struct Branch {
	BranchJson // mut:
}
