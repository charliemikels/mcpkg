module main

struct BranchJson {}
struct Branch {
	BranchJson
	// mut:
}
