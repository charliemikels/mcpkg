module main
// main.v is currently for testing purposes and should be phased out once mcpkg-cli exists.

fn main() {
	println('hello again.')
}
